* C:\Users\Zulfiqar\Desktop\supply\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sun Dec 12 21:08:18 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END

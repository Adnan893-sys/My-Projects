* C:\Users\Zulfiqar\Desktop\supply\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Sun Dec 12 22:03:08 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
